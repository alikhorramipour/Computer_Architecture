----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:53:11 05/15/2019 
-- Design Name: 
-- Module Name:    cc - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;
entity CPU8BIT2 is
port ( data: out std_logic_vector(7 downto 0);
	adress: out std_logic_vector(5 downto 0);
	oe: out std_logic;
	we: out std_logic; -- Asynchronous memory interface
	rst: in std_logic;
	clk: in std_logic);
end;
architecture CPU_ARCH of CPU8BIT2 is
signal akku: std_logic_vector(8 downto 0); -- akku(8) is carry !
signal adreg: std_logic_vector(4 downto 0);
signal pc: std_logic_vector(4 downto 0);
signal clock: std_logic;
signal states: std_logic_vector(2 downto 0);
type memory is array(32 downto 0) of std_logic_vector(7 downto 0);
	begin
	Process(clock,rst)
		begin
		If (rst = '0') then
			adreg <= (others => '0'); -- start execution at memory location 0
			states <= "000";
			akku <= (others => '0');
			pc <= (others => '0');
		elsIf rising_edge(clk) then
		-- PC / Adress path
			If (states = "000") then
				pc <= adreg + 1;
				adreg <= my_Rom(To_integer(unsigned(pc)))(4 downto 0);
			else
				adreg <= pc;
			end If;
			-- ALU / Data Path
			Case states is
			when "001" => akku <= ("0" & akku(7 downto 0)) - ("0" & my_Rom(To_integer(unsigned(adreg ))));
			when "010" => akku <= ("0" & akku(7 downto 0)) + ("0" & my_Rom(To_integer(unsigned(adreg )))); -- add
			when "011" => akku(7 downto 0) <= akku(7 downto 0) nor my_Rom(To_integer(unsigned(adreg ))); -- nor
			when "100" => akku(8) <= '0'; -- branch not taken, clear carry
			when "101" => akku <= (others => '0');
			when "110" => akku <= ("0" & akku(7 downto 0)) xor ("0" & my_Rom(To_integer(unsigned(adreg ))));
			when "111" => akku <= ("0" & akku(7 downto 0)) and ("0" & my_Rom(To_integer(unsigned(adreg ))));
			when others => null; -- instr. fetch, jcc taken (000), sta (001)
		end Case;
		-- State machine
		If (states /= "000") then states <= "000"; -- fetch next opcode
		else states <=  not my_Rom(To_integer(unsigned(pc)))(7 downto 5); -- execute instruction
		end If;
		end If;
		end Process;
		-- output
		adress <= '0'&adreg;
		data <= akku(7 downto 0);
		oe <= '1' when (clk='1' or states = "001" or rst='0' or states = "101") else '0';
		-- no memory access during reset and state "101" (branch not taken)
		we <= '1' when (clk='1' or states /= "001" or rst='0') else '0';
end CPU_ARCH;