--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:06:31 05/29/2019
-- Design Name:   
-- Module Name:   D:/407 - 426/J11/tbPipelined.vhd
-- Project Name:  J11
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Pipelined
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tbPipelined IS
END tbPipelined;
 
ARCHITECTURE behavior OF tbPipelined IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Pipelined
    PORT(
         clock : IN  std_logic;
			rst : IN  std_logic;
         a : IN  std_logic_vector(1 downto 0);
         b : IN  std_logic_vector(1 downto 0);
         c : IN  std_logic_vector(1 downto 0);
         data : IN  std_logic_vector(1 downto 0);
         result : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clock : std_logic := '0';
   signal a : std_logic_vector(1 downto 0) := (others => '0');
   signal b : std_logic_vector(1 downto 0) := (others => '0');
   signal c : std_logic_vector(1 downto 0) := (others => '0');
   signal data : std_logic_vector(1 downto 0) := (others => '0');
	signal rst : std_logic := '0';
 	
	--Outputs
   signal result : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clock_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Pipelined PORT MAP (
          clock => clock,
          a => a,
          b => b,
          c => c,
          data => data,
          result => result,
			 rst => rst
        );

   -- Clock process definitions
   clock_process :process
   begin
		clock <= '0';
		wait for clock_period/2;
		clock <= '1';
		wait for clock_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		rst <= '0';
		a <= "10";
		b <= "01";
		c <= "11";
		data <= "10";
		
      wait for 100 ns;	

      wait for clock_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
